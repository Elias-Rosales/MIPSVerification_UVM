parameter DMEMORY_WIDTH = 100;